netcdf ini_hydro {

dimensions:
	xi_rho = 130 ;
	xi_u = 129 ;
	xi_v = 130 ;
	eta_rho = 130 ;
	eta_u = 130 ;
	eta_v = 129 ;
	s_rho = 20 ;
	s_w = 21 ;
	tracer = 2 ;
	time = UNLIMITED ; // (0 currently)

variables:
	char spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:option_T = "spherical" ;
		spherical:option_F = "Cartesian" ;
	double ocean_time(time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 0000-01-01 00:00:00" ;
		ocean_time:calendar = "360.0 days in every year" ;
		ocean_time:field = "time, scalar, series" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
		theta_s:units = "nondimensional" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
		theta_b:units = "nondimensional" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:units = "nondimensional" ;
		s_rho:valid_min = 0. ;
		s_rho:valid_max = -1. ;
                s_rho:formula_terms = "s: s_rho eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:units = "nondimensional" ;
		s_w:valid_min = 0. ;
		s_w:valid_max = -1. ;
                s_w:standard_name = "ocean_s_coordinate" ;
                s_w:formula_terms = "s: s_w eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:units = "nondimensional" ;
		Cs_r:valid_min = 0. ;
		Cs_r:valid_max = -1. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:units = "nondimensional" ;
		Cs_w:valid_min = 0. ;
		Cs_w:valid_max = -1. ;
		Cs_w:field = "Cs_w, scalar" ;
	double zeta(time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:field = "free-surface, scalar, series" ;
		zeta:time = "ocean_time" ;
	double ubar(time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:field = "ubar-velocity, scalar, series" ;
		ubar:time = "ocean_time" ;
	double vbar(time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:field = "vbar-velocity, scalar, series" ;
		vbar:time = "ocean_time" ;
	double u(time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:field = "u-velocity, scalar, series" ;
		u:time = "ocean_time" ;
	double v(time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:field = "v-velocity, scalar, series" ;
		v:time = "ocean_time" ;
	double temp(time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:field = "temperature, scalar, series" ;
		temp:time = "ocean_time" ;
	double salt(time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:units = "PSU" ;
		salt:field = "salinity, scalar, series" ;
		salt:time = "ocean_time" ;

// global attributes:
		:type = "INITIALIZATION file" ;
		:title = "Levitus One-degree Annual Climatology (1994) - DAMEE # 4" ;
		:out_file = "damee4_levfeb.nc" ;
		:grd_file = "damee4_grid_a.nc" ;
		:history = "Version 4.0  , Tuesday - March 14, 2000 - 5:04:02 PM" ;

}
