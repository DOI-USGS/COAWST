netcdf ini_sed {

dimensions:
	xi_rho = 102 ;
	xi_u = 101 ;
	xi_v = 102 ;
	xi_psi = 101 ;
	eta_rho = 22 ;
	eta_u = 22 ;
	eta_v = 21 ;
	eta_psi = 21 ;
	s_rho = 8 ;
	s_w = 9 ;
	tracer = 3 ;
	Nbed = 1 ;
	time = UNLIMITED ; // (0 currently)

variables:
	char spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:option_T = "spherical" ;
		spherical:option_F = "Cartesian" ;
	double ocean_time(time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 0000-01-01 00:00:00" ;
		ocean_time:calendar = "365.25 days in every year" ;
		ocean_time:field = "time, scalar, series" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
		theta_s:units = "nondimensional" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
		theta_b:units = "nondimensional" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:units = "nondimensional" ;
		s_rho:valid_min = 0. ;
		s_rho:valid_max = -1. ;
                s_rho:formula_terms = "s: s_rho eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:units = "nondimensional" ;
		s_w:valid_min = 0. ;
		s_w:valid_max = -1. ;
                s_w:standard_name = "ocean_s_coordinate" ;
                s_w:formula_terms = "s: s_w eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:units = "nondimensional" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:units = "nondimensional" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
		Cs_w:field = "Cs_w, scalar" ;
	float zeta(time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:field = "free-surface, scalar, series" ;
	float ubar(time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:field = "ubar-velocity, scalar, series" ;
	float vbar(time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:field = "vbar-velocity, scalar, series" ;
	float u(time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
		u:field = "u-velocity, scalar, series" ;
	float v(time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
		v:field = "v-velocity, scalar, series" ;
	float w(time, s_w, eta_rho, xi_rho) ;
		w:long_name = "vertical momentum component" ;
		w:units = "meter second-1" ;
		w:time = "ocean_time" ;
		w:field = "w-velocity, scalar, series" ;
	float omega(time, s_w, eta_rho, xi_rho) ;
		omega:long_name = "S-coordinate vertical momentum component" ;
		omega:units = "meter3 second-1" ;
		omega:time = "ocean_time" ;
		omega:field = "omega, scalar, series" ;
	float temp(time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:time = "ocean_time" ;
		temp:field = "temperature, scalar, series" ;
	float salt(time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:units = "PSU" ;
		salt:time = "ocean_time" ;
		salt:field = "salinity, scalar, series" ;
	float mud_01(time, s_rho, eta_rho, xi_rho) ;
		mud_01:long_name = "suspended cohesive sediment, size class 01" ;
		mud_01:size_class = " 1.0000E-02 millimeter" ;
		mud_01:units = "milligram liter-1" ;
		mud_01:time = "ocean_time" ;
		mud_01:field = "mud_01, scalar, series" ;
	float mudfrac_01(time, Nbed, eta_rho, xi_rho) ;
		mudfrac_01:long_name = "cohesive sediment fraction, size class 01" ;
		mudfrac_01:size_class = " 1.0000E-02 millimeter" ;
		mudfrac_01:units = "nondimensional" ;
		mudfrac_01:time = "ocean_time" ;
		mudfrac_01:field = "mudfrac_01, scalar, series" ;
	float mudmass_01(time, Nbed, eta_rho, xi_rho) ;
		mudmass_01:long_name = "cohesive sediment mass, size class 01" ;
		mudmass_01:size_class = " 1.0000E-02 millimeter" ;
		mudmass_01:units = "kilogram meter-2" ;
		mudmass_01:time = "ocean_time" ;
		mudmass_01:field = "mudmass_01, scalar, series" ;
	float bed_thickness(time, Nbed, eta_rho, xi_rho) ;
		bed_thickness:long_name = "sediment layer thickness" ;
		bed_thickness:units = "meter" ;
		bed_thickness:time = "ocean_time" ;
		bed_thickness:field = "bed_thickness, scalar, series" ;
	float bed_age(time, Nbed, eta_rho, xi_rho) ;
		bed_age:long_name = "sediment layer age" ;
		bed_age:units = "day" ;
		bed_age:time = "ocean_time" ;
		bed_age:field = "bed_age, scalar, series" ;
	float bed_porosity(time, Nbed, eta_rho, xi_rho) ;
		bed_porosity:long_name = "sediment layer porosity" ;
		bed_porosity:units = "nondimensional" ;
		bed_porosity:time = "ocean_time" ;
		bed_porosity:field = "bed_porosity, scalar, series" ;
	float grain_size(time, eta_rho, xi_rho) ;
		grain_size:long_name = "sediment median grain diameter size" ;
		grain_size:units = "meter" ;
		grain_size:time = "ocean_time" ;
		grain_size:field = "grain_size, scalar, series" ;
	float grain_density(time, eta_rho, xi_rho) ;
		grain_density:long_name = "sediment medina grain density" ;
		grain_density:units = "kilogram meter3" ;
		grain_density:time = "ocean_time" ;
		grain_density:field = "grain_density, scalar, series" ;
	float settling_vel(time, eta_rho, xi_rho) ;
		settling_vel:long_name = "sediment median grain settling velocity" ;
		settling_vel:units = "meter second-1" ;
		settling_vel:time = "ocean_time" ;
		settling_vel:field = "settling_vel, scalar, series" ;
	float erosion_stress(time, eta_rho, xi_rho) ;
		erosion_stress:long_name = "sediment median critical erosion stress" ;
		erosion_stress:units = "meter2 second-2" ;
		erosion_stress:time = "ocean_time" ;
		erosion_stress:field = "erosion_stress, scalar, series" ;
	float bed_wave_amp(time, eta_rho, xi_rho) ;
		bed_wave_amp:long_name = "bed wave excursion amplitude" ;
		bed_wave_amp:units = "meter" ;
		bed_wave_amp:time = "ocean_time" ;
		bed_wave_amp:field = "bed_wave_amp, scalar, series" ;

// global attributes:
		:type = "ROMS INITIAL file" ;
		:title = "ROMS Initial fiels for Hydrodynamics and Sediment" ;
		:grd_file = "roms_grd.nc" ;

}
