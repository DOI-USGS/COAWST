netcdf bry_unlimit {

dimensions:
	xi_rho = 66 ;
	eta_rho = 194 ;
	xi_u = 65 ;
	eta_u = 194 ;
	xi_v = 66 ;
	eta_v = 193 ;
	s_rho = 30 ;
	bry_time = UNLIMITED ; // (0 currently)

variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "open boundary conditions time" ;
		bry_time:units = "days since 0000-01-01 00:00:00" ;
		bry_time:field = "bry_time, scalar, series" ;
	float zeta_west(bry_time, eta_rho) ;
		zeta_west:long_name = "free-surface western boundary condition" ;
		zeta_west:units = "meter" ;
		zeta_west:field = "zeta_west, scalar, series" ;
		zeta_west:time = "bry_time" ;
	float zeta_east(bry_time, eta_rho) ;
		zeta_east:long_name = "free-surface eastern boundary condition" ;
		zeta_east:units = "meter" ;
		zeta_east:field = "zeta_east, scalar, series" ;
		zeta_east:time = "bry_time" ;
	float zeta_south(bry_time, xi_rho) ;
		zeta_south:long_name = "free-surface southern boundary condition" ;
		zeta_south:units = "meter" ;
		zeta_south:field = "zeta_south, scalar, series" ;
		zeta_south:time = "bry_time" ;
	float zeta_north(bry_time, xi_rho) ;
		zeta_north:long_name = "free-surface northern boundary condition" ;
		zeta_north:units = "meter" ;
		zeta_north:field = "zeta_north, scalar, series" ;
		zeta_north:time = "bry_time" ;
	float ubar_west(bry_time, eta_u) ;
		ubar_west:long_name = "2D u-momentum western boundary condition" ;
		ubar_west:units = "meter second-1" ;
		ubar_west:field = "ubar_west, scalar, series" ;
		ubar_west:time = "bry_time" ;
	float ubar_east(bry_time, eta_u) ;
		ubar_east:long_name = "2D u-momentum eastern boundary condition" ;
		ubar_east:units = "meter second-1" ;
		ubar_east:field = "ubar_east, scalar, series" ;
		ubar_east:time = "bry_time" ;
	float ubar_south(bry_time, xi_u) ;
		ubar_south:long_name = "2D u-momentum southern boundary condition" ;
		ubar_south:units = "meter second-1" ;
		ubar_south:field = "ubar_south, scalar, series" ;
		ubar_south:time = "bry_time" ;
	float ubar_north(bry_time, xi_u) ;
		ubar_north:long_name = "2D u-momentum northern boundary condition" ;
		ubar_north:units = "meter second-1" ;
		ubar_north:field = "ubar_north, scalar, series" ;
		ubar_north:time = "bry_time" ;
	float vbar_west(bry_time, eta_v) ;
		vbar_west:long_name = "2D v-momentum western boundary condition" ;
		vbar_west:units = "meter second-1" ;
		vbar_west:field = "vbar_west, scalar, series" ;
		vbar_west:time = "bry_time" ;
	float vbar_east(bry_time, eta_v) ;
		vbar_east:long_name = "2D v-momentum eastern boundary condition" ;
		vbar_east:units = "meter second-1" ;
		vbar_east:field = "vbar_east, scalar, series" ;
		vbar_east:time = "bry_time" ;
	float vbar_south(bry_time, xi_v) ;
		vbar_south:long_name = "2D v-momentum southern boundary condition" ;
		vbar_south:units = "meter second-1" ;
		vbar_south:field = "vbar_south, scalar, series" ;
		vbar_south:time = "bry_time" ;
	float vbar_north(bry_time, xi_v) ;
		vbar_north:long_name = "2D v-momentum northern boundary condition" ;
		vbar_north:units = "meter second-1" ;
		vbar_north:field = "vbar_north, scalar, series" ;
		vbar_north:time = "bry_time" ;
	float u_west(bry_time, s_rho, eta_u) ;
		u_west:long_name = "3D u-momentum western boundary condition" ;
		u_west:units = "meter second-1" ;
		u_west:field = "u_west, scalar, series" ;
		u_west:time = "bry_time" ;
	float u_east(bry_time, s_rho, eta_u) ;
		u_east:long_name = "3D u-momentum eastern boundary condition" ;
		u_east:units = "meter second-1" ;
		u_east:field = "u_east, scalar, series" ;
		u_east:time = "bry_time" ;
	float u_south(bry_time, s_rho, xi_u) ;
		u_south:long_name = "3D u-momentum southern boundary condition" ;
		u_south:units = "meter second-1" ;
		u_south:field = "u_south, scalar, series" ;
		u_south:time = "bry_time" ;
	float u_north(bry_time, s_rho, xi_u) ;
		u_north:long_name = "3D u-momentum northern boundary condition" ;
		u_north:units = "meter second-1" ;
		u_north:field = "u_north, scalar, series" ;
		u_north:time = "bry_time" ;
	float v_west(bry_time, s_rho, eta_v) ;
		v_west:long_name = "3D v-momentum western boundary condition" ;
		v_west:units = "meter second-1" ;
		v_west:field = "v_west, scalar, series" ;
		v_west:time = "bry_time" ;
	float v_east(bry_time, s_rho, eta_v) ;
		v_east:long_name = "3D v-momentum eastern boundary condition" ;
		v_east:units = "meter second-1" ;
		v_east:field = "v_east, scalar, series" ;
		v_east:time = "bry_time" ;
	float v_south(bry_time, s_rho, xi_v) ;
		v_south:long_name = "3D v-momentum southern boundary condition" ;
		v_south:units = "meter second-1" ;
		v_south:field = "v_south, scalar, series" ;
		v_south:time = "bry_time" ;
	float v_north(bry_time, s_rho, xi_v) ;
		v_north:long_name = "3D v-momentum northern boundary condition" ;
		v_north:units = "meter second-1" ;
		v_north:field = "v_north, scalar, series" ;
		v_north:time = "bry_time" ;
	float temp_west(bry_time, s_rho, eta_rho) ;
		temp_west:long_name = "potential temperature western boundary condition" ;
		temp_west:units = "Celsius" ;
		temp_west:field = "temp_west, scalar, series" ;
		temp_west:time = "bry_time" ;
	float temp_east(bry_time, s_rho, eta_rho) ;
		temp_east:long_name = "potential temperature eastern boundary condition" ;
		temp_east:units = "Celsius" ;
		temp_east:field = "temp_east, scalar, series" ;
		temp_east:time = "bry_time" ;
	float temp_south(bry_time, s_rho, xi_rho) ;
		temp_south:long_name = "potential temperature southern boundary condition" ;
		temp_south:units = "Celsius" ;
		temp_south:field = "temp_south, scalar, series" ;
		temp_south:time = "bry_time" ;
	float temp_north(bry_time, s_rho, xi_rho) ;
		temp_north:long_name = "potential temperature northern boundary condition" ;
		temp_north:units = "Celsius" ;
		temp_north:field = "temp_north, scalar, series" ;
		temp_north:time = "bry_time" ;
	float salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity western boundary condition" ;
		salt_west:units = "PSU" ;
		salt_west:field = "salt_west, scalar, series" ;
		salt_west:time = "bry_time" ;
	float salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity eastern boundary condition" ;
		salt_east:units = "PSU" ;
		salt_east:field = "salt_east, scalar, series" ;
		salt_east:time = "bry_time" ;
	float salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity southern boundary condition" ;
		salt_south:units = "PSU" ;
		salt_south:field = "salt_south, scalar, series" ;
		salt_south:time = "bry_time" ;
	float salt_north(bry_time, s_rho, xi_rho) ;
		salt_north:long_name = "salinity northern boundary condition" ;
		salt_north:units = "PSU" ;
		salt_north:field = "salt_north, scalar, series" ;
		salt_north:time = "bry_time" ;

// global attributes:
		:type = "BOUNDARY FORCING file" ;
		:title = "Northeast North American (NENA) Shelf Model" ;
		:grd_file = "roms_nena_grid_2.nc" ;
		:history = "BOUNDARY file, 1.0  , 27-Mar-2002 13:11:22" ;

}
