netcdf clm_ts {

dimensions:
	xi_rho = 130 ;
	xi_u = 129 ;
	xi_v = 130 ;
	eta_rho = 130 ;
	eta_u = 130 ;
	eta_v = 129 ;
	s_rho = 20 ;
	s_w = 21 ;
	tracer = 2 ;
	temp_time = 12 ;
	salt_time = 12 ;

variables:
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
		theta_s:units = "nondimensional" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
		theta_b:units = "nondimensional" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:units = "nondimensional" ;
		s_rho:valid_min = 0. ;
		s_rho:valid_max = -1. ;
                s_rho:formula_terms = "s: s_rho eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:units = "nondimensional" ;
		s_w:valid_min = 0. ;
		s_w:valid_max = -1. ;
                s_w:standard_name = "ocean_s_coordinate" ;
                s_w:formula_terms = "s: s_w eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:units = "nondimensional" ;
		Cs_r:valid_min = 0. ;
		Cs_r:valid_max = -1. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:units = "nondimensional" ;
		Cs_w:valid_min = 0. ;
		Cs_w:valid_max = -1. ;
		Cs_w:field = "Cs_w, scalar" ;
	double temp_time(temp_time) ;
		temp_time:long_name = "time for potential temperature" ;
		temp_time:units = "day" ;
		temp_time:field = "temp_time, scalar, series" ;
		temp_time:cycle_length = 360. ;
	double salt_time(salt_time) ;
		salt_time:long_name = "time for salinity" ;
		salt_time:units = "day" ;
		salt_time:field = "salt_time, scalar, series" ;
		salt_time:cycle_length = 360. ;
	float temp(temp_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:field = "temperature, scalar, series" ;
		temp:time = "temp_time" ;
	float salt(salt_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:units = "PSU" ;
		salt:field = "salinity, scalar, series" ;
		salt:time = "salt_time" ;

// global attributes:
		:type = "CLIMATOLOGY file" ;
		:title = "Levitus One-Degree Monthly T-S Climatology (1994) - DAMEE #4" ;
		:out_file = "damee4_Lclm.nc" ;
		:grd_file = "damee4_grid_a.nc" ;
		:history = "Version 4.0  , Tuesday - March 21, 2000 - 4:47:16 PM" ;

}
