netcdf adriatic1_frc {
dimensions:
	xi_rho = 42 ;
	eta_rho = 142 ;
	xi_u = 41 ;
	eta_u = 142 ;
	xi_v = 42 ;
	eta_v = 141 ;
        zeta_time = 12;
	v2d_time = 12 ;
	v3d_time = 12 ;
	temp_time = 12 ;
	salt_time = 12 ;
variables:
	double zeta_time(zeta_time) ;
		zeta_time:long_name = "free-surface time" ;
		zeta_time:units = "days since 0000-01-01 00:00:00" ;
		zeta_time:field = "zeta_time, scalar, series" ;
		zeta_time:cycle_length = 360. ;
	double v2d_time(v2d_time) ;
		v2d_time:long_name = "2D momentum time" ;
		v2d_time:units = "days since 0000-01-01 00:00:00" ;
		v2d_time:field = "v2d_time, scalar, series" ;
		v2d_time:cycle_length = 360. ;
	double v3d_time(v3d_time) ;
		v3d_time:long_name = "3D momentum time" ;
		v3d_time:units = "days since 0000-01-01 00:00:00" ;
		v3d_time:field = "v3d_time, scalar, series" ;
		v3d_time:cycle_length = 360. ;
	double temp_time(temp_time) ;
		temp_time:long_name = "potential temperature time" ;
		temp_time:units = "days since 0000-01-01 00:00:00" ;
		temp_time:field = "temp_time, scalar, series" ;
		temp_time:cycle_length = 360. ;
	double salt_time(salt_time) ;
		salt_time:long_name = "surface net heat flux time" ;
		salt_time:units = "days since 0000-01-01 00:00:00" ;
		salt_time:field = "salt_time, scalar, series" ;
		salt_time:cycle_length = 360. ;
	float zeta_west(zeta_time, eta_rho) ;
		zeta_west:long_name = "free-surface western boundary condition" ;
		zeta_west:units = "meter" ;
		zeta_west:field = "zeta_west, scalar, series" ;
		zeta_west:time = "zeta_time" ;
	float zeta_east(zeta_time, eta_rho) ;
		zeta_east:long_name = "free-surface eastern boundary condition" ;
		zeta_east:units = "meter" ;
		zeta_east:field = "zeta_east, scalar, series" ;
		zeta_east:time = "zeta_time" ;
	float zeta_south(zeta_time, xi_rho) ;
		zeta_south:long_name = "free-surface southern boundary condition" ;
		zeta_south:units = "meter" ;
		zeta_south:field = "zeta_south, scalar, series" ;
		zeta_south:time = "zeta_time" ;
	float zeta_north(zeta_time, xi_rho) ;
		zeta_north:long_name = "free-surface northern boundary condition" ;
		zeta_north:units = "meter" ;
		zeta_north:field = "zeta_north, scalar, series" ;
		zeta_north:time = "zeta_time" ;
	float ubar_west(v2d_time, eta_u) ;
		ubar_west:long_name = "2D u-momentum western boundary condition" ;
		ubar_west:units = "meter second-1" ;
		ubar_west:field = "ubar_west, scalar, series" ;
		ubar_west:time = "v2d_time" ;
	float ubar_east(v2d_time, eta_u) ;
		ubar_east:long_name = "2D u-momentum eastern boundary condition" ;
		ubar_east:units = "meter second-1" ;
		ubar_east:field = "ubar_east, scalar, series" ;
		ubar_east:time = "v2d_time" ;
	float ubar_south(v2d_time, xi_u) ;
		ubar_south:long_name = "2D u-momentum southern boundary condition" ;
		ubar_south:units = "meter second-1" ;
		ubar_south:field = "ubar_south, scalar, series" ;
		ubar_south:time = "v2d_time" ;
	float ubar_north(v2d_time, xi_u) ;
		ubar_north:long_name = "2D u-momentum northern boundary condition" ;
		ubar_north:units = "meter second-1" ;
		ubar_north:field = "ubar_north, scalar, series" ;
		ubar_north:time = "v2d_time" ;
	float vbar_west(v2d_time, eta_v) ;
		vbar_west:long_name = "2D v-momentum western boundary condition" ;
		vbar_west:units = "meter second-1" ;
		vbar_west:field = "vbar_west, scalar, series" ;
		vbar_west:time = "v2d_time" ;
	float vbar_east(v2d_time, eta_v) ;
		vbar_east:long_name = "2D v-momentum eastern boundary condition" ;
		vbar_east:units = "meter second-1" ;
		vbar_east:field = "vbar_east, scalar, series" ;
		vbar_east:time = "v2d_time" ;
	float vbar_south(v2d_time, xi_v) ;
		vbar_south:long_name = "2D v-momentum southern boundary condition" ;
		vbar_south:units = "meter second-1" ;
		vbar_south:field = "vbar_south, scalar, series" ;
		vbar_south:time = "v2d_time" ;
	float vbar_north(v2d_time, xi_v) ;
		vbar_north:long_name = "2D v-momentum northern boundary condition" ;
		vbar_north:units = "meter second-1" ;
		vbar_north:field = "vbar_north, scalar, series" ;
		vbar_north:time = "v2d_time" ;
	float u_west(v3d_time, s_rho, eta_u) ;
		u_west:long_name = "3D u-momentum western boundary condition" ;
		u_west:units = "meter second-1" ;
		u_west:field = "u_west, scalar, series" ;
		u_west:time = "v3d_time" ;
	float u_east(v3d_time, s_rho, eta_u) ;
		u_east:long_name = "3D u-momentum eastern boundary condition" ;
		u_east:units = "meter second-1" ;
		u_east:field = "u_east, scalar, series" ;
		u_east:time = "v3d_time" ;
	float u_south(v3d_time, s_rho, xi_u) ;
		u_south:long_name = "3D u-momentum southern boundary condition" ;
		u_south:units = "meter second-1" ;
		u_south:field = "u_south, scalar, series" ;
		u_south:time = "v3d_time" ;
	float u_north(v3d_time, s_rho, xi_u) ;
		u_north:long_name = "3D u-momentum northern boundary condition" ;
		u_north:units = "meter second-1" ;
		u_north:field = "u_north, scalar, series" ;
		u_north:time = "v3d_time" ;
	float v_west(v3d_time, s_rho, eta_v) ;
		v_west:long_name = "3D v-momentum western boundary condition" ;
		v_west:units = "meter second-1" ;
		v_west:field = "v_west, scalar, series" ;
		v_west:time = "v3d_time" ;
	float v_east(v3d_time, s_rho, eta_v) ;
		v_east:long_name = "3D v-momentum eastern boundary condition" ;
		v_east:units = "meter second-1" ;
		v_east:field = "v_east, scalar, series" ;
		v_east:time = "v3d_time" ;
	float v_south(v3d_time, s_rho, xi_v) ;
		v_south:long_name = "3D v-momentum southern boundary condition" ;
		v_south:units = "meter second-1" ;
		v_south:field = "v_south, scalar, series" ;
		v_south:time = "v3d_time" ;
	float v_north(v3d_time, s_rho, xi_v) ;
		v_north:long_name = "3D v-momentum northern boundary condition" ;
		v_north:units = "meter second-1" ;
		v_north:field = "v_north, scalar, series" ;
		v_north:time = "v3d_time" ;
	float temp_west(temp_time, s_rho, eta_rho) ;
		temp_west:long_name = "potential temperature western boundary condition" ;
		temp_west:units = "Celsius" ;
		temp_west:field = "temp_west, scalar, series" ;
		temp_west:time = "temp_time" ;
	float temp_east(temp_time, s_rho, eta_rho) ;
		temp_east:long_name = "potential temperature eastern boundary condition" ;
		temp_east:units = "Celsius" ;
		temp_east:field = "temp_east, scalar, series" ;
		temp_east:time = "temp_time" ;
	float temp_south(temp_time, s_rho, xi_rho) ;
		temp_south:long_name = "potential temperature southern boundary condition" ;
		temp_south:units = "Celsius" ;
		temp_south:field = "temp_south, scalar, series" ;
		temp_south:time = "temp_time" ;
	float temp_north(temp_time, s_rho, xi_rho) ;
		temp_north:long_name = "potential temperature northern boundary condition" ;
		temp_north:units = "Celsius" ;
		temp_north:field = "temp_north, scalar, series" ;
		temp_north:time = "temp_time" ;
	float salt_west(salt_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity western boundary condition" ;
		salt_west:units = "PSU" ;
		salt_west:field = "salt_west, scalar, series" ;
		salt_west:time = "salt_time" ;
	float salt_east(salt_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity eastern boundary condition" ;
		salt_east:units = "PSU" ;
		salt_east:field = "salt_east, scalar, series" ;
		salt_east:time = "salt_time" ;
	float salt_south(salt_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity southern boundary condition" ;
		salt_south:units = "PSU" ;
		salt_south:field = "salt_south, scalar, series" ;
		salt_south:time = "salt_time" ;
	float salt_north(salt_time, s_rho, xi_rho) ;
		salt_north:long_name = "salinity northern boundary condition" ;
		salt_north:units = "PSU" ;
		salt_north:field = "salt_north, scalar, series" ;
		salt_north:time = "salt_time" ;

// global attributes:
		:title = "Adriatic Boundary Forcing, Grid # 1" ;
		:history = "BOUNDARY file, 4.0  , Tuesday - April 2, 2002 - 6:29:46 PM" ;
		:type = "BOUNDARY FORCING file" ;
		:out_file = "adriatic1_frc.nc" ;
		:grd_file = "adriatic1_grd.nc" ;

data:

 zeta_time = 15, 45, 75, 105, 135, 165, 195, 225, 255, 285, 315, 345 ;

 v2d_time = 15, 45, 75, 105, 135, 165, 195, 225, 255, 285, 315, 345 ;

 v3d_time = 15, 45, 75, 105, 135, 165, 195, 225, 255, 285, 315, 345 ;

 temp_time = 15, 45, 75, 105, 135, 165, 195, 225, 255, 285, 315, 345 ;

 salt_time = 15, 45, 75, 105, 135, 165, 195, 225, 255, 285, 315, 345 ;

}
