netcdf grd_spherical {

dimensions:
	xi_psi = 110 ;
	xi_rho = 111 ;
	xi_u = 110 ;
	xi_v = 111 ;
	eta_psi = 240 ;
	eta_rho = 241 ;
	eta_u = 241 ;
	eta_v = 240 ;
	bath = UNLIMITED ; // (0 currently)

variables:
	char spherical ;
		spherical:long_name = "Grid type logical switch" ;
		spherical:option_T = "spherical" ;
		spherical:option_F = "Cartesian" ;
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	double hraw(bath, eta_rho, xi_rho) ;
		hraw:long_name = "Working bathymetry at RHO-points" ;
		hraw:units = "meter" ;
		hraw:field = "bath, scalar" ;
	double h(eta_rho, xi_rho) ;
		h:long_name = "Final bathymetry at RHO-points" ;
		h:units = "meter" ;
		h:field = "bath, scalar" ;
	double f(eta_rho, xi_rho) ;
		f:long_name = "Coriolis parameter at RHO-points" ;
		f:units = "second-1" ;
		f:field = "Coriolis, scalar" ;
	double pm(eta_rho, xi_rho) ;
		pm:long_name = "curvilinear coordinate metric in XI" ;
		pm:units = "meter-1" ;
		pm:field = "pm, scalar" ;
	double pn(eta_rho, xi_rho) ;
		pn:long_name = "curvilinear coordinate metric in ETA" ;
		pn:units = "meter-1" ;
		pn:field = "pn, scalar" ;
	double dndx(eta_rho, xi_rho) ;
		dndx:long_name = "xi derivative of inverse metric factor pn" ;
		dndx:units = "meter" ;
		dndx:field = "dndx, scalar" ;
	double dmde(eta_rho, xi_rho) ;
		dmde:long_name = "eta derivative of inverse metric factor pm" ;
		dmde:units = "meter" ;
		dmde:field = "dmde, scalar" ;
	double x_rho(eta_rho, xi_rho) ;
		x_rho:long_name = "x location of RHO-points" ;
		x_rho:units = "meter" ;
	double y_rho(eta_rho, xi_rho) ;
		y_rho:long_name = "y location of RHO-points" ;
		y_rho:units = "meter" ;
	double x_psi(eta_psi, xi_psi) ;
		x_psi:long_name = "x location of PSI-points" ;
		x_psi:units = "meter" ;
	double y_psi(eta_psi, xi_psi) ;
		y_psi:long_name = "y location of PSI-points" ;
		y_psi:units = "meter" ;
	double x_u(eta_u, xi_u) ;
		x_u:long_name = "x location of U-points" ;
		x_u:units = "meter" ;
	double y_u(eta_u, xi_u) ;
		y_u:long_name = "y location of U-points" ;
		y_u:units = "meter" ;
	double x_v(eta_v, xi_v) ;
		x_v:long_name = "x location of V-points" ;
		x_v:units = "meter" ;
	double y_v(eta_v, xi_v) ;
		y_v:long_name = "y location of V-points" ;
		y_v:units = "meter" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
	double lat_psi(eta_psi, xi_psi) ;
		lat_psi:long_name = "latitude of PSI-points" ;
		lat_psi:units = "degree_north" ;
	double lon_psi(eta_psi, xi_psi) ;
		lon_psi:long_name = "longitude of PSI-points" ;
		lon_psi:units = "degree_east" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
        double angle(eta_rho, xi_rho) ;
                angle:long_name = "angle between XI-axis and EAST" ;
                angle:units = "radians" ;
                angle:field = "angle, scalar" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:option_0 = "land" ;
		mask_rho:option_1 = "water" ;
		mask_rho:_FillValue = 1. ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:option_0 = "land" ;
		mask_u:option_1 = "water" ;
		mask_u:_FillValue = 1. ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:option_0 = "land" ;
		mask_v:option_1 = "water" ;
		mask_v:_FillValue = 1. ;
	double mask_psi(eta_psi, xi_psi) ;
		mask_psi:long_name = "mask on PSI-points" ;
		mask_psi:option_0 = "land" ;
		mask_psi:option_1 = "water" ;
		mask_psi:_FillValue = 1. ;

// global attributes:
		:type = "ROMS GRID file" ;
		:title = "NJB grid for LEO-15" ;

}
